module scope
module chk